library verilog;
use verilog.vl_types.all;
entity testIIR is
end testIIR;
