library verilog;
use verilog.vl_types.all;
entity testmul is
end testmul;
