library verilog;
use verilog.vl_types.all;
entity testIIR_look_ahead_pipe is
end testIIR_look_ahead_pipe;
