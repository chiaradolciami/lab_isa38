library verilog;
use verilog.vl_types.all;
entity test_fpmult is
end test_fpmult;
